library verilog;
use verilog.vl_types.all;
entity score_to_bcd_vlg_vec_tst is
end score_to_bcd_vlg_vec_tst;
