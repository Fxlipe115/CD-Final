library verilog;
use verilog.vl_types.all;
entity clock_count_vlg_vec_tst is
end clock_count_vlg_vec_tst;
