library verilog;
use verilog.vl_types.all;
entity sequence_vlg_vec_tst is
end sequence_vlg_vec_tst;
