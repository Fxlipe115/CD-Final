library verilog;
use verilog.vl_types.all;
entity genius_vlg_vec_tst is
end genius_vlg_vec_tst;
